//Subject:     CO project 2 - Sign extend
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      
//----------------------------------------------
//Date:        
//----------------------------------------------
//Description: 
//--------------------------------------------------------------------------------
//add zero or one  to the offset's left side by this offset  pos or neg [15]
`timescale 1ns/1ps
module Sign_Extend(
    data_i,
    data_o
    );
               
//I/O ports
input   [16-1:0] data_i;
output  [32-1:0] data_o;

//Internal Signals
reg     [32-1:0] data_o;

//Sign extended
always @(data_i) begin
	data_o[15:0] <= data_i[15:0];
	//positive
	if (data_i[15]==0) 
		data_o[31:16] <= 16'b0;
	//negative
	else 
		data_o[31:16] <= ~(16'b0);
end
endmodule      
     